`timescale 1ns / 1ps
module Mux2to1_4bit (
    input [3:0] A, B,  // ????????? ? ????
    input S,           // ?????? ?????? (0: A, 1: B)
    input E,           // ?????? ????????? (0: ????, 1: ???????)
    output [3:0] Y     // ????? ? ????
);
    // ?????? ???? ?? ????? ????
    assign Y = (E == 1'b1) ? 4'bzzzz :  // ??? E=1? ????? High-Z
               (S == 1'b0) ? A : B;     // ??? E=0? ?????? A ?? B ?????? S
endmodule